----------------------------------------------------------------------------------
-- TECHNICAL UNIVERSITY OF CRETE
-- NICK KYPARISSAS
--
-- CREATE DATE: JUNE 2018
-- MODULE NAME: TOP LEVEL MODULE
-- PROJECT NAME: A Parallel Framework for Simulating Cellular Automata on FPGA Logic
-- XILINX OPEN HARDWARE 2018 ENTRY
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TOP_LEVEL IS
	GENERIC ( 	GRID_X				: INTEGER := 1920; -- NUMBER OF CELLS IN A LINE 
				GRID_Y				: INTEGER := 1080; -- NUMBER OF LINES
				CELL_SIZE  			: INTEGER := 4;--8; 
				-- CELL SIZE IN BITS
				-- CELL_SIZE = 4 => 2^4 = 16 STATES
				-- CELL_SIZE = 8 => 2^8 = 256 STATES 
				BURST_SIZE 			: INTEGER := 128; -- NUMBER OF BITS
				NUMBER_OF_BURSTS_PER_LINE 	: INTEGER := 60;--120;
				-- CELL_SIZE = 4 => NUMBER_OF_BURSTS_PER_LINE = GRID_X * CELL_SIZE / BURST_SIZE = 60
				-- CELL_SIZE = 8 => NUMBER_OF_BURSTS_PER_LINE = GRID_X * CELL_SIZE / BURST_SIZE = 120
        		NEIGHBORHOOD_SIZE  	: INTEGER := 21; -- NEIGHBORHOOD SIZE MUST BE AN ODD NUMBER >= 3
        		-- SPEED: EVERY N FRAMES => NEW GENERATION
        		-- FOR EXAMPLE, OUR GRAPHICS HERE RUN AT 60 FPS. 
        		-- IF SPEED = 60: A NEW GENERATION WILL BE CALCULATED EVERY 1 SEC
        		MEMORY_ADDR_WIDTH	: INTEGER := 27 -- NUMBER OF BITS
	);
    PORT ( 	
		CLK					: IN STD_LOGIC;	-- EXTERNAL CLOCK
		RST 				: IN STD_LOGIC;
		-- GRAPHICS SIGNALS --
		HS          : OUT STD_LOGIC;
		VS          : OUT STD_LOGIC;
		R           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		G           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		B           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		-- MEMORY SIGNALS --
		DDR2_DQ     : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		DDR2_DQS_P  : INOUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		DDR2_DQS_N  : INOUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		DDR2_ADDR   : OUT   STD_LOGIC_VECTOR(12 DOWNTO 0);
		DDR2_BA     : OUT   STD_LOGIC_VECTOR(2 DOWNTO 0);
		DDR2_RAS_N  : OUT   STD_LOGIC;
		DDR2_CAS_N  : OUT   STD_LOGIC;
		DDR2_WE_N   : OUT   STD_LOGIC;
		DDR2_CK_P   : OUT   STD_LOGIC_VECTOR(0 DOWNTO 0);
		DDR2_CK_N   : OUT   STD_LOGIC_VECTOR(0 DOWNTO 0);
		--ddr2_cs_n	: OUT   STD_LOGIC_VECTOR(0 DOWNTO 0);
		DDR2_CKE    : OUT   STD_LOGIC_VECTOR(0 DOWNTO 0);
		DDR2_DM     : OUT   STD_LOGIC_VECTOR(1 DOWNTO 0);
		DDR2_ODT    : OUT   STD_LOGIC_VECTOR(0 DOWNTO 0);
		-- UART SIGNALS --
		UART_RX 	: IN  STD_LOGIC;
		-- SPEED CONTROL
		SPEED_UP    : IN STD_LOGIC;
		SPEED_DOWN  : IN STD_LOGIC;
		-- OPERATIONAL INDICATORS [LEDS] --
		UART_OP				: OUT STD_LOGIC;
        GRAPHICS_MEM_ACCESS_OP : OUT STD_LOGIC;
        CA_ENGINE_MEM_ACCESS_OP : OUT STD_LOGIC;
		INIT_COMPLETE_OP 	: OUT STD_LOGIC;
		APP_RDY_OP : OUT STD_LOGIC;
		APP_WDF_RDY_OP : OUT STD_LOGIC
	);
END TOP_LEVEL;

ARCHITECTURE BEHAVIORAL OF TOP_LEVEL IS
	
	-- CLOCKING WIZARD SIGNALS --
	SIGNAL CLK325_SIGNAL, CLK200_SIGNAL, CLK148_SIGNAL : STD_LOGIC;
	
	-- UART SIGNALS --
	SIGNAL UART_RX_DATA : STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL UART_RX_DATA_RDY, UART_FRAME_ERROR : STD_LOGIC := '0';
	
	-- UART FIFO SIGNALS --
	SIGNAL INIT_UART_FIFO_DATA_SIGNAL : STD_LOGIC_VECTOR(127 DOWNTO 0) := (OTHERS => '0');
	SIGNAL INIT_UART_FIFO_READ_EN_SIGNAL : STD_LOGIC := '0';
	SIGNAL INIT_UART_FIFO_EMPTY_SIGNAL : STD_LOGIC := '1';
	
	-- INITIALIZATION FIFO HANDLER SIGNALS -- 
	SIGNAL APP_EN_INIT_SIGNAL, APP_WDF_END_INIT_SIGNAL, APP_WDF_WREN_INIT_SIGNAL : STD_LOGIC := '0';
    SIGNAL INIT_COMPLETE_SIGNAL : STD_LOGIC := '0';
	SIGNAL APP_CMD_INIT_SIGNAL : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
	SIGNAL APP_WDF_DATA_INIT_SIGNAL : STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL APP_ADDR_INIT_SIGNAL  	: STD_LOGIC_VECTOR(MEMORY_ADDR_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
	
	-- GRAPHICS BUFFER SIGNALS --
	SIGNAL APP_EN_GRAPHICS_SIGNAL, GRAPHICS_FIFO_FULL_SIGNAL, GRAPHICS_MEM_EN_SIGNAL : STD_LOGIC := '0';
	SIGNAL APP_CMD_GRAPHICS_SIGNAL : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
	SIGNAL APP_ADDR_GRAPHICS_SIGNAL  : STD_LOGIC_VECTOR(MEMORY_ADDR_WIDTH-1 DOWNTO 0) := (OTHERS => '0');	
	SIGNAL GRAPHICS_DATA_SIGNAL	: STD_LOGIC_VECTOR(127 DOWNTO 0) := (OTHERS => '0');
	
	-- DATAPATH FEEDER SIGNALS --
	SIGNAL NEIGHBORHOOD_DATA_SIGNAL : STD_LOGIC_VECTOR((NEIGHBORHOOD_SIZE*CELL_SIZE)-1 DOWNTO 0) := (OTHERS  => '0');
	
	-- CA ENGINE SIGNALS --
	SIGNAL LINE_BUFFER_DATA_VALID : STD_LOGIC := '0';
	SIGNAL CA_ENGINE_DATA_OUT_SIGNAL : STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL CA_ENGINE_FIFO_WRITE_EN_SIGNAL, CA_ENGINE_FIFO_EMPTY_SIGNAL : STD_LOGIC := '0';
        
	-- WRITE-BACK SIGNALS -- 
	SIGNAL WRITE_BACK_FIFO_DATA_SIGNAL : STD_LOGIC_VECTOR(127 DOWNTO 0) := (OTHERS => '0');
	SIGNAL APP_EN_WRITE_BACK_SIGNAL, APP_WDF_END_WRITE_BACK_SIGNAL, APP_WDF_WREN_WRITE_BACK_SIGNAL, WRITE_BACK_FIFO_READY_SIGNAL, WRITE_BACK_FIFO_READ_EN_SIGNAL : STD_LOGIC := '0';
	SIGNAL APP_CMD_WRITE_BACK_SIGNAL : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
	SIGNAL APP_WDF_DATA_WRITE_BACK_SIGNAL : STD_LOGIC_VECTOR(127 DOWNTO 0) := (OTHERS => '0');
	SIGNAL APP_ADDR_WRITE_BACK_SIGNAL : STD_LOGIC_VECTOR(MEMORY_ADDR_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
	 
	-- MEMORY ACCESS CONTROL --
	SIGNAL GRAPHICS_ACCESS_REQ_SIGNAL, GRAPHICS_ACCESS_GRANTED_SIGNAL, GRAPHICS_NEW_FRAME_REQ_SIGNAL, WRITE_BACK_ACCESS_GRANTED_SIGNAL : STD_LOGIC := '0'; -- PIPELINING_SIGNAL VERSION ABOVE (WE DONT CARE IF THEY ARE LATE - INDEPENDENTLY STALL SOMETHING IRRELEVANT TO THEIR SOURCE)
	SIGNAL APP_CMD_SELECT_SIGNAL : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0'); -- 00: INIT, 01: READING BUFFER, 10: WRITING BUFFER, 11: GRAPHICS BUFFER
	SIGNAL APP_WRITE_SELECT_SIGNAL : STD_LOGIC := '0'; -- 0: INIT, 1: WRITING BUFFER	
	
	-- MEMORY INTERFACE GENERATOR/SOLUTION (MIG/S) SIGNALS --
	SIGNAL UI_CLK_SIGNAL : STD_LOGIC;
	SIGNAL APP_RDY_SIGNAL, APP_RD_DATA_VALID_SIGNAL, APP_WDF_RDY_SIGNAL, APP_EN_SIGNAL, APP_WDF_END_SIGNAL, APP_WDF_WREN_SIGNAL :  STD_LOGIC := '0';
	SIGNAL APP_CMD_SIGNAL : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
	SIGNAL APP_WDF_DATA_SIGNAL, APP_RD_DATA_SIGNAL	: STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAl APP_ADDR_SIGNAL	: STD_LOGIC_VECTOR(MEMORY_ADDR_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
	
	-- MISC SIGNALS
	SIGNAL SPEED : INTEGER RANGE 0 TO 30 := 30;
	
	
	-- COMPONENTS
	COMPONENT mig_7series_0 
	port (
		ddr2_dq : inout std_logic_vector(15 downto 0);
		ddr2_dqs_p : inout std_logic_vector(1 downto 0);
		ddr2_dqs_n : inout std_logic_vector(1 downto 0);
		ddr2_addr  : out   std_logic_vector(12 downto 0);
		ddr2_ba : out   std_logic_vector(2 downto 0);
		ddr2_ras_n : out std_logic;
		ddr2_cas_n : out std_logic;
		ddr2_we_n : out std_logic;
		ddr2_ck_p : out std_logic_vector(0 downto 0);
		ddr2_ck_n : out std_logic_vector(0 downto 0);
		ddr2_cke : out std_logic_vector(0 downto 0);
		ddr2_dm : out std_logic_vector(1 downto 0);
		ddr2_odt : out std_logic_vector(0 downto 0);
		app_addr : in std_logic_vector(26 downto 0);
		app_cmd : in std_logic_vector(2 downto 0);
		app_en : in std_logic;
		app_wdf_data : in std_logic_vector(127 downto 0);
		app_wdf_end : in std_logic;
		app_wdf_mask : in std_logic_vector(15 downto 0);
		app_wdf_wren : in std_logic;
		app_rd_data : out std_logic_vector(127 downto 0);
		app_rd_data_end : out std_logic;
		app_rd_data_valid : out std_logic;
		app_rdy : out std_logic;
		app_wdf_rdy : out std_logic;
		app_sr_req : in std_logic;
		app_ref_req : in std_logic;
		app_zq_req : in std_logic;
		app_sr_active : out std_logic;
		app_ref_ack : out std_logic;
		app_zq_ack: out std_logic;
		ui_clk : out std_logic;
		ui_clk_sync_rst : out std_logic;
		init_calib_complete : out std_logic;
		-- System Clock Ports
		sys_clk_i : in std_logic;
		-- Reference Clock Ports
		clk_ref_i : in std_logic;
		sys_rst : in std_logic
	);
	END COMPONENT;
	
	COMPONENT clk_wiz_0
	PORT ( 
		clk_out1 	: OUT STD_LOGIC; -- 200 MHz
		clk_out2 	: OUT STD_LOGIC; -- 325 MHz
		reset 		: IN STD_LOGIC;
		locked      : OUT STD_LOGIC;
		clk_in 		: IN STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT clk_wiz_1 
	PORT (
		clk_out1 	: OUT STD_LOGIC; -- 148.5 MHz
		reset 		: IN STD_LOGIC;
		clk_in 		: IN STD_LOGIC
	);
	END COMPONENT;
	
	COMPONENT GRAPHICS_FIFO
        PORT (
		rst : IN STD_LOGIC;
		wr_clk : IN STD_LOGIC;
		rd_clk : IN STD_LOGIC;
		din : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		wr_en : IN STD_LOGIC;
		rd_en : IN STD_LOGIC;
		dout : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		full : OUT STD_LOGIC;
		empty : OUT STD_LOGIC
	);
    END COMPONENT;	
	BEGIN
	
	CLOCKING_WIZARD: clk_wiz_0  
	PORT MAP(
		clk_out1 => CLK200_SIGNAL, -- 200 MHz, DDR reference CLK (required: +- 200 MHz)
		clk_out2 => CLK325_SIGNAL, -- 325 MHz (required: +- 324.9 MHz)
		reset => RST, 
		clk_in => CLK
	);
	
	CLOCKING_WIZARD_GRAPHICS: clk_wiz_1 
	PORT MAP(
		clk_out1 => CLK148_SIGNAL, -- 148 MHz, for graphics (required: +- 148.5 MHz)
		reset => RST,  
		clk_in => CLK
	);

    GRAPHICS_BUFFER: GRAPHICS_FIFO
    PORT MAP (
        rst => RST,
        wr_clk => UI_CLK_SIGNAL, 
        rd_clk => CLK148_SIGNAL,
        din => APP_RD_DATA_SIGNAL,
        wr_en => APP_RD_DATA_VALID_SIGNAL,
        rd_en => GRAPHICS_MEM_EN_SIGNAL,
        dout => GRAPHICS_DATA_SIGNAL,
        full => GRAPHICS_FIFO_FULL_SIGNAL
	);
    
    MIG_CONTROLLER: mig_7series_0 
	PORT MAP(
		DDR2_DQ => DDR2_DQ,   
		DDR2_DQS_P => DDR2_DQS_P,
		DDR2_DQS_N => DDR2_DQS_N,
		DDR2_ADDR => DDR2_ADDR, 
		DDR2_BA => DDR2_BA,   
		DDR2_RAS_N => DDR2_RAS_N,
		DDR2_CAS_N => DDR2_CAS_N,
		DDR2_WE_N => DDR2_WE_N,
		DDR2_CK_P => DDR2_CK_P,
		DDR2_CK_N => DDR2_CK_N,
		DDR2_CKE => DDR2_CKE,
		DDR2_DM => DDR2_DM, 
		DDR2_ODT => DDR2_ODT,
		APP_ADDR => APP_ADDR_SIGNAL,
		APP_CMD => APP_CMD_SIGNAL, 
		APP_EN => APP_EN_SIGNAL,
		APP_WDF_DATA => APP_WDF_DATA_SIGNAL,
		APP_WDF_END => APP_WDF_END_SIGNAL,
		APP_WDF_MASK => (OTHERS => '0'),
		APP_WDF_WREN => APP_WDF_WREN_SIGNAL,
		APP_RD_DATA => APP_RD_DATA_SIGNAL,
		APP_RD_DATA_VALID => APP_RD_DATA_VALID_SIGNAL,
		APP_RDY => APP_RDY_SIGNAL,
		APP_WDF_RDY => APP_WDF_RDY_SIGNAL,
		APP_SR_REQ => '0',
		APP_REF_REQ => '0',
		APP_ZQ_REQ => '0',         
		UI_CLK => UI_CLK_SIGNAL,  
		SYS_CLK_I => CLK325_SIGNAL, -- 325 MHz (required: +- 324.9 MHz)
		clk_ref_i => CLK200_SIGNAL, -- 196.3 MHz (required: +- 200 MHz)
		SYS_RST => RST
	);

	UART_CONTROLLER: ENTITY WORK.UART 
    PORT MAP(
        CLK         => CLK,
        RST         => RST,
        -- UART INTERFACE
        UART_RXD    => UART_RX,
        -- USER DATA INPUT INTERFACE
        DATA_IN  => "00000000",
        DATA_SEND => '0', 
        -- USER DATA OUTPUT INTERFACE
        DATA_OUT => UART_RX_DATA,
        DATA_VLD  => UART_RX_DATA_RDY,
        FRAME_ERROR => UART_FRAME_ERROR 
    );
    
    INIT_UART_FIFO: ENTITY WORK.FIFO_8_128
    PORT MAP (
        -- WRITE PORT
        din => UART_RX_DATA,
        wr_en => UART_RX_DATA_RDY,
        -- READ PORT
        rd_en => INIT_UART_FIFO_READ_EN_SIGNAL,
        dout => INIT_UART_FIFO_DATA_SIGNAL,
        empty => INIT_UART_FIFO_EMPTY_SIGNAL,
        ------------
        rst => RST,
        wr_clk => CLK,
        rd_clk => UI_CLK_SIGNAL
    );
	
	MEMORY_INITIALIZER: ENTITY WORK.MEMORY_INITIALIZER
	GENERIC MAP (
		CELL_SIZE => CELL_SIZE,
		BURST_SIZE => BURST_SIZE,
		NUMBER_OF_BURSTS_PER_LINE => NUMBER_OF_BURSTS_PER_LINE,
		GRID_Y => GRID_Y,
		MEMORY_ADDR_WIDTH => MEMORY_ADDR_WIDTH
	)
    PORT MAP (
		CLK => UI_CLK_SIGNAL, -- 81.25MHZ FROM DDR'S UI_CLK
		RST => RST,
		-- CONTROL SIGNALS --
		INIT_COMPLETE => INIT_COMPLETE_SIGNAL,
		-- FIFO HANDLING SIGNALS --
		FIFO_DATA => INIT_UART_FIFO_DATA_SIGNAL,
		FIFO_READ_EN => INIT_UART_FIFO_READ_EN_SIGNAL,
		FIFO_EMPTY => INIT_UART_FIFO_EMPTY_SIGNAL,
		-- MEMORY SIGNALS --- 
		APP_RDY => APP_RDY_SIGNAL,
		APP_WDF_RDY => APP_WDF_RDY_SIGNAL,
		APP_EN => APP_EN_INIT_SIGNAL,
		APP_CMD => APP_CMD_INIT_SIGNAL, 
		APP_WDF_DATA => APP_WDF_DATA_INIT_SIGNAL,
		APP_WDF_END => APP_WDF_END_INIT_SIGNAL,
		APP_WDF_WREN => APP_WDF_WREN_INIT_SIGNAL,
		APP_ADDR => APP_ADDR_INIT_SIGNAL
	);
	
	MEMORY_ACCESS_ARBITRATOR: ENTITY WORK.MEMORY_ACCESS_ARBITRATOR
    PORT MAP( 	
		CLK	=> UI_CLK_SIGNAL, --CLK1_SIGNAL
		RST => RST,
		-- INIT SIGNALS --
		INIT_COMPLETE => INIT_COMPLETE_SIGNAL, 
		-- GRAPHICS SIGNALS	--
		GRAPHICS_REQ => GRAPHICS_ACCESS_REQ_SIGNAL,
		GRAPHICS_NEW_FRAME_REQ => GRAPHICS_NEW_FRAME_REQ_SIGNAL,
		GRAPHICS_ACCESS_GRANTED	=> GRAPHICS_ACCESS_GRANTED_SIGNAL, 
		-- WRITING BUFFER SIGNALS --
		WRITE_BACK_ACCESS_GRANTED => WRITE_BACK_ACCESS_GRANTED_SIGNAL,
		-- DDR SIGNALS --
		APP_CMD_SELECT => APP_CMD_SELECT_SIGNAL, 
		APP_WRITE_SELECT => APP_WRITE_SELECT_SIGNAL			
	);
	
	MEMORY_CMD_MUX: ENTITY WORK.DDR_CMD_MUX 
	PORT MAP(
		APP_ADDR_INIT => APP_ADDR_INIT_SIGNAL,
		APP_CMD_INIT => APP_CMD_INIT_SIGNAL,
		APP_EN_INIT => APP_EN_INIT_SIGNAL,
		APP_ADDR_WRITE => APP_ADDR_WRITE_BACK_SIGNAL,
		APP_CMD_WRITE => APP_CMD_WRITE_BACK_SIGNAL,
		APP_EN_WRITE => APP_EN_WRITE_BACK_SIGNAL,		
		APP_ADDR_GRAPHICS => APP_ADDR_GRAPHICS_SIGNAL,		
		APP_CMD_GRAPHICS => APP_CMD_GRAPHICS_SIGNAL,
		APP_EN_GRAPHICS	=> APP_EN_GRAPHICS_SIGNAL,
		SEL => APP_CMD_SELECT_SIGNAL, 
		APP_ADDR => APP_ADDR_SIGNAL,
		APP_CMD	=> APP_CMD_SIGNAL,
		APP_EN	=> APP_EN_SIGNAL
	);
		
	MEMORY_WRITE_MUX: ENTITY WORK.DDR_WRITE_MUX 
	PORT MAP(
        APP_WDF_DATA_INIT => APP_WDF_DATA_INIT_SIGNAL,
		APP_WDF_END_INIT => APP_WDF_END_INIT_SIGNAL,
		APP_WDF_WREN_INIT => APP_WDF_WREN_INIT_SIGNAL,
		APP_WDF_DATA_WRITE => APP_WDF_DATA_WRITE_BACK_SIGNAL,
		APP_WDF_END_WRITE  => APP_WDF_END_WRITE_BACK_SIGNAL,
		APP_WDF_WREN_WRITE	 => APP_WDF_WREN_WRITE_BACK_SIGNAL,
        SEL => APP_WRITE_SELECT_SIGNAL,
		APP_WDF_DATA => APP_WDF_DATA_SIGNAL,
		APP_WDF_END	=> APP_WDF_END_SIGNAL,
		APP_WDF_WREN => APP_WDF_WREN_SIGNAL
	);
	
	GRAPHICS_FEEDER: ENTITY WORK.GRAPHICS_FEEDER 
    GENERIC MAP ( 	
				MEMORY_ADDRESS_WIDTH => MEMORY_ADDR_WIDTH,
				GRID_Y => GRID_Y,
				NUMBER_OF_BURSTS_PER_LINE => NUMBER_OF_BURSTS_PER_LINE
	)
    PORT MAP ( 	
		CLK	=> UI_CLK_SIGNAL,
		RST => RST,
		-- CONTROL SIGNALS --
		MEM_ACCESS_GRANTED	=> GRAPHICS_ACCESS_GRANTED_SIGNAL,
		SPEED => SPEED,		
		-- MEMORY SIGNALS --
		APP_RDY => APP_RDY_SIGNAL,
		APP_ADDR => APP_ADDR_GRAPHICS_SIGNAL,
		APP_EN => APP_EN_GRAPHICS_SIGNAL,
		APP_CMD => APP_CMD_GRAPHICS_SIGNAL
	);
    
	GRAPHICS_CONTROLLER: ENTITY WORK.GRAPHICS_CTRL
	GENERIC MAP ( 	
	   COLOR_BITS => CELL_SIZE
	)
	PORT MAP( 
		CLK => CLK148_SIGNAL,
		RST => RST,
		MEM_DATA => GRAPHICS_DATA_SIGNAL,
		MEM_EN => GRAPHICS_MEM_EN_SIGNAL,
		HS => HS,
        VS => VS,
		MEM_ACCESS_REQUEST => GRAPHICS_ACCESS_REQ_SIGNAL,
		NEW_FRAME_LINE_REQUEST => GRAPHICS_NEW_FRAME_REQ_SIGNAL,
        R => R,
        G => G,
        B => B
	);
	
	CA_ENGINE_WRITE_BACK: ENTITY WORK.WRITE_BACK
	GENERIC MAP ( 	
			MEMORY_ADDRESS_WIDTH => MEMORY_ADDR_WIDTH,
			NUMBER_OF_ROWS	=> GRID_Y,
			NEIGHBORHOOD_SIZE => NEIGHBORHOOD_SIZE,
			NUMBER_OF_BURSTS_PER_LINE => NUMBER_OF_BURSTS_PER_LINE,
			BURST_SIZE => BURST_SIZE
	)
	PORT MAP(
		CLK	=> UI_CLK_SIGNAL,
		RST => RST,
		-- CONTROL SIGNALS --
		MEM_ACCESS_GRANTED => WRITE_BACK_ACCESS_GRANTED_SIGNAL,
		-- FIFO SIGNALS
		FIFO_DATA => WRITE_BACK_FIFO_DATA_SIGNAL,
		FIFO_READ_EN => WRITE_BACK_FIFO_READ_EN_SIGNAL,
		FIFO_READY => WRITE_BACK_FIFO_READY_SIGNAL,
		--
		SPEED => SPEED,
		-- MEMORY SIGNALS --
		APP_RDY => APP_RDY_SIGNAL,
		APP_WDF_RDY => APP_WDF_RDY_SIGNAL,
		APP_EN => APP_EN_WRITE_BACK_SIGNAL,
		APP_CMD => APP_CMD_WRITE_BACK_SIGNAL,
		APP_WDF_DATA => APP_WDF_DATA_WRITE_BACK_SIGNAL,
		APP_WDF_END => APP_WDF_END_WRITE_BACK_SIGNAL,
		APP_WDF_WREN => APP_WDF_WREN_WRITE_BACK_SIGNAL,
		APP_ADDR => APP_ADDR_WRITE_BACK_SIGNAL
	);
	

	WRITE_BACK_FIFO_4: IF (CELL_SIZE = 4) GENERATE
		WRITE_BACK_FIFO: ENTITY WORK.FIFO_4_128
	    PORT MAP (
	        -- WRITE PORT
	        din => CA_ENGINE_DATA_OUT_SIGNAL,
	        wr_en => CA_ENGINE_FIFO_WRITE_EN_SIGNAL,
	        -- READ PORT
	        rd_en => WRITE_BACK_FIFO_READ_EN_SIGNAL,
	        dout => WRITE_BACK_FIFO_DATA_SIGNAL,
	        empty => CA_ENGINE_FIFO_EMPTY_SIGNAL, 
	        ------------
	        rst => RST,
	        wr_clk => CLK200_SIGNAL,
	        rd_clk => UI_CLK_SIGNAL
	    );
	END GENERATE;
	
	WRITE_BACK_FIFO_8:	IF (CELL_SIZE = 8) GENERATE
		WRITE_BACK_FIFO_8: ENTITY WORK.FIFO_8_128
	    PORT MAP (
	        -- WRITE PORT
	        din => CA_ENGINE_DATA_OUT_SIGNAL,
	        wr_en => CA_ENGINE_FIFO_WRITE_EN_SIGNAL,
	        -- READ PORT
	        rd_en => WRITE_BACK_FIFO_READ_EN_SIGNAL,
	        dout => WRITE_BACK_FIFO_DATA_SIGNAL,
	        empty => CA_ENGINE_FIFO_EMPTY_SIGNAL, 
	        ------------
	        rst => RST,
	        wr_clk => CLK200_SIGNAL,
	        rd_clk => UI_CLK_SIGNAL
	    );
    END GENERATE;
    
    WRITE_BACK_FIFO_READY_SIGNAL <=  NOT CA_ENGINE_FIFO_EMPTY_SIGNAL;
 
	GRID_LINES_BUFFER: ENTITY WORK.GRID_LINES_BUFFER
	GENERIC MAP (
        CELL_SIZE => CELL_SIZE,		
		BURST_SIZE => BURST_SIZE,
		GRID_X => GRID_X,
		GRID_Y => GRID_Y,
		NUMBER_OF_BURSTS_PER_LINE => NUMBER_OF_BURSTS_PER_LINE,
        NEIGHBORHOOD_SIZE => NEIGHBORHOOD_SIZE
    ) 
	PORT MAP(
        CLK_200 => CLK200_SIGNAL,
		UI_CLK => UI_CLK_SIGNAL,
        RST => RST,
		WRITE_EN => APP_RD_DATA_VALID_SIGNAL,
		MEMORY_ACCESS_GRANTED => GRAPHICS_ACCESS_GRANTED_SIGNAL,
        DATA_IN => APP_RD_DATA_SIGNAL,
        DATA_OUT => NEIGHBORHOOD_DATA_SIGNAL,
        DATA_OUT_VALID => LINE_BUFFER_DATA_VALID
        );
	
    CA_ENGINE: ENTITY WORK.CA_ENGINE
    GENERIC MAP (
            CELL_SIZE => CELL_SIZE,
            NEIGHBORHOOD_SIZE => NEIGHBORHOOD_SIZE
    )
    PORT MAP ( 
    	CLK => CLK200_SIGNAL,
    	RST => RST,
    	
    	READ_EN => LINE_BUFFER_DATA_VALID,
    	DATA_IN => NEIGHBORHOOD_DATA_SIGNAL,
    	
    	DATA_OUT => CA_ENGINE_DATA_OUT_SIGNAL,
        DATA_OUT_VALID => CA_ENGINE_FIFO_WRITE_EN_SIGNAL    	
    );
    
    SPEED_CONTROLLER: PROCESS
    BEGIN
    
        WAIT UNTIL RISING_EDGE(UI_CLK_SIGNAL);
        
        IF RST = '1' THEN
            SPEED <= 30;
        ELSE
            IF SPEED_DOWN = '1' AND SPEED < 30 THEN
                SPEED <= SPEED + 10;            
            ELSIF SPEED_UP = '1' AND SPEED > 0 THEN
                SPEED <= SPEED - 10; 
            ELSE
                SPEED <= SPEED;       
            END IF;
        END IF;
        
    END PROCESS;
    
    -- OPERATIONAL INDICATORS [LEDS] --
	UART_OP	<= (UART_RX_DATA(3) OR UART_RX_DATA(2) OR UART_RX_DATA(1) OR UART_RX_DATA(0)) AND (NOT INIT_COMPLETE_SIGNAL); -- VALID, INCOMING DATA
	INIT_COMPLETE_OP <= INIT_COMPLETE_SIGNAL;
	--
	GRAPHICS_MEM_ACCESS_OP <= GRAPHICS_ACCESS_GRANTED_SIGNAL;
    CA_ENGINE_MEM_ACCESS_OP <= WRITE_BACK_ACCESS_GRANTED_SIGNAL; 
    --  
	APP_RDY_OP <= APP_RDY_SIGNAL;
	APP_WDF_RDY_OP <= APP_WDF_RDY_SIGNAL;
	
	END BEHAVIORAL;