----------------------------------------------------------------------------------
-- TECHNICAL UNIVERSITY OF CRETE
-- NICK KYPARISSAS
--
-- CREATE DATE: JUNE 2018
-- MODULE: Ca Engine implementing the "HODGEPODGE MACHINE" rule
-- PROJECT NAME: A Parallel Framework for Simulating Cellular Automata on FPGA Logic
-- XILINX OPEN HARDWARE 2018 ENTRY
----------------------------------------------------------------------------------

-- YOU CANT USE THIS AS IS: EVERY TIME THE NEIGHBORHOOD SIZE CHANGES, 
-- THE ADDERS BINARY TREE MIGHT REQUIRE CHANGES AS WELL. 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CA_ENGINE IS
	GENERIC (
        CELL_SIZE   	: INTEGER := 8; -- HOW MANY BITS PER CELL - WIDTH MUST BE DIVIDED BY CELL SIZE
        NEIGHBORHOOD_SIZE : INTEGER := 21);  -- OUTPUT DATA DEPTH IN CELLS - ARRAY DEPTH
        -- FOR EXAMPLE: IF WIDTH = 7 CELLS, CELL SIZE = 4 BITS AND DEPTH = 7 CELLS, THEN 
        -- DATA IN = 32 CELLS = 32*4 BITS = 128 BITS (IN MY APPLICATION: THIS WAS THE MEMORY BURST SIZE)
        -- DATA OUT = 7 CELLS = 7*4 BITS = 28 BITS
    PORT  ( 
    	CLK : IN STD_LOGIC;
    	RST : IN STD_LOGIC;
    	
    	READ_EN : IN STD_LOGIC;
    	DATA_IN : IN STD_LOGIC_VECTOR((NEIGHBORHOOD_SIZE*CELL_SIZE)-1 DOWNTO 0);
    	
    	DATA_OUT : OUT STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
        DATA_OUT_VALID : OUT STD_LOGIC
    	
    );
END CA_ENGINE;

ARCHITECTURE BEHAVIORAL OF CA_ENGINE IS

-- PIPELINED NEIGHBORHOOD
type NEIGHBORHOOD_ARRAY is array (NEIGHBORHOOD_SIZE-1 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 255; -- 256 STATES
SIGNAL NEIGHBORHOOD_CELL, NEIGHBORHOOD_REPLICA : NEIGHBORHOOD_ARRAY := (OTHERS => (OTHERS => 0));

-- EACH ARRAY CELL MUST BE LARGE ENOUGH FOR NEIGHBORHOOD_CELL*NEIGHBORHOOD_WEIGHT
type CATEGORIZED_NEIGHBORHOOD_ARRAY is array (NEIGHBORHOOD_SIZE-1 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 1;
SIGNAL INFECTED_CELL, ILL_CELL : CATEGORIZED_NEIGHBORHOOD_ARRAY := (OTHERS => (OTHERS => 0));

-- YOU NEED TO ADJUST THIS SIGNAL ACCORDING TO THE DEPTH OF YOUR RULE'S PIPELINE 
SIGNAL DATA_VALID_SIGNAL : STD_LOGIC_VECTOR( ((NEIGHBORHOOD_SIZE-1)/2)+12 DOWNTO 0) := (OTHERS => '0');

-- CUSTOM RULE SIGNALS
-- TREE OF SUMS FOR THE STATES SUM
type SUM_LAYER_0_TYPE is array ((NEIGHBORHOOD_SIZE-1)/2 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 93000;
SIGNAL SUM_LAYER_0 : SUM_LAYER_0_TYPE;
type SUM_LAYER_1_TYPE is array ((NEIGHBORHOOD_SIZE-1)/4 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 93000;
SIGNAL SUM_LAYER_1 : SUM_LAYER_1_TYPE;
type SUM_LAYER_2_TYPE is array (2 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 93000;
SIGNAL SUM_LAYER_2 : SUM_LAYER_2_TYPE;
type SUM_LAYER_3_TYPE is array (1 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 93000;
SIGNAL SUM_LAYER_3 : SUM_LAYER_3_TYPE;		
type SUM_TYPE is array (NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 93000;
SIGNAL SUM : SUM_TYPE;	
type COLUMN_SUM_LAYER_0_TYPE is array ((NEIGHBORHOOD_SIZE-1)/2 downto 0) of integer range 0 to 93000;
SIGNAL COLUMN_SUM_LAYER_0 : COLUMN_SUM_LAYER_0_TYPE;
type COLUMN_SUM_LAYER_1_TYPE is array ((NEIGHBORHOOD_SIZE-1)/4 downto 0) of integer range 0 to 93000;
SIGNAL COLUMN_SUM_LAYER_1 : COLUMN_SUM_LAYER_1_TYPE;
type COLUMN_SUM_LAYER_2_TYPE is array (2 downto 0) of integer range 0 to 93000;
SIGNAL COLUMN_SUM_LAYER_2 : COLUMN_SUM_LAYER_2_TYPE;
type COLUMN_SUM_LAYER_3_TYPE is array (1 downto 0) of integer range 0 to 93000;
SIGNAL COLUMN_SUM_LAYER_3 : COLUMN_SUM_LAYER_3_TYPE;		
SIGNAL TOTAL_SUM : integer range 0 to 93000;	

-- TREE OF SUMS FOR THE TOTAL NUMBER OF INFECTED CELLS
type INFECTED_SUM_LAYER_0_TYPE is array ((NEIGHBORHOOD_SIZE-1)/2 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_SUM_LAYER_0 : INFECTED_SUM_LAYER_0_TYPE;
type INFECTED_SUM_LAYER_1_TYPE is array ((NEIGHBORHOOD_SIZE-1)/4 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_SUM_LAYER_1 : INFECTED_SUM_LAYER_1_TYPE;
type INFECTED_SUM_LAYER_2_TYPE is array (2 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_SUM_LAYER_2 : INFECTED_SUM_LAYER_2_TYPE;
type INFECTED_SUM_LAYER_3_TYPE is array (1 downto 0, NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_SUM_LAYER_3 : INFECTED_SUM_LAYER_3_TYPE;		
type INFECTED_SUM_TYPE is array (NEIGHBORHOOD_SIZE-1 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_SUM : INFECTED_SUM_TYPE;	
type INFECTED_COLUMN_SUM_LAYER_0_TYPE is array ((NEIGHBORHOOD_SIZE-1)/2 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_COLUMN_SUM_LAYER_0 : INFECTED_COLUMN_SUM_LAYER_0_TYPE;
type INFECTED_COLUMN_SUM_LAYER_1_TYPE is array ((NEIGHBORHOOD_SIZE-1)/4 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_COLUMN_SUM_LAYER_1 : INFECTED_COLUMN_SUM_LAYER_1_TYPE;
type INFECTED_COLUMN_SUM_LAYER_2_TYPE is array (2 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_COLUMN_SUM_LAYER_2 : INFECTED_COLUMN_SUM_LAYER_2_TYPE;
type INFECTED_COLUMN_SUM_LAYER_3_TYPE is array (1 downto 0) of integer range 0 to 511;
SIGNAL INFECTED_COLUMN_SUM_LAYER_3 : INFECTED_COLUMN_SUM_LAYER_3_TYPE;		
SIGNAL INFECTED_TOTAL_SUM : integer range 0 to 511;	

TYPE CURRENT_CELL_PIPELINE is array (222 downto 0) of integer range 0 to 255;
SIGNAL CURRENT_CELL : CURRENT_CELL_PIPELINE := (OTHERS => 0);
	
SIGNAL SUM_DIVIDED : STD_LOGIC_VECTOR(16 DOWNTO 0);	
	
BEGIN
     
	PROCESS 
	BEGIN
		
		WAIT UNTIL RISING_EDGE(CLK);	
		
		IF RST = '1' THEN
			DATA_VALID_SIGNAL <= (OTHERS => '0');
		END IF;
		
		-- PIPELINING NEIGHBORHOOD ----------------------------------
        FOR I IN NEIGHBORHOOD_SIZE-1 DOWNTO 1 LOOP
            FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 0 LOOP
                NEIGHBORHOOD_CELL(I, J) <= NEIGHBORHOOD_CELL(I-1, J);
            END LOOP;
        END LOOP;
        
        FOR I IN NEIGHBORHOOD_SIZE-1 DOWNTO 0 LOOP
            NEIGHBORHOOD_CELL(0, I) <= TO_INTEGER(UNSIGNED(DATA_IN((I*CELL_SIZE)+CELL_SIZE-1 DOWNTO I*CELL_SIZE)));
        END LOOP;
        
        -- SETTING UP THE 3 DIFFERENT ADDER TREES
        FOR I IN NEIGHBORHOOD_SIZE-1 DOWNTO 0 LOOP
            FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 0 LOOP
                NEIGHBORHOOD_REPLICA(I, J) <= NEIGHBORHOOD_CELL(I, J);
            	IF NEIGHBORHOOD_CELL(I, J) > 0 THEN
                	INFECTED_CELL(I, J) <= 1;
           	 	ELSE
            		INFECTED_CELL(I, J) <= 0;
            	END IF;                
            END LOOP;
        END LOOP;
        
        FOR I IN 10 DOWNTO 1 LOOP
        	CURRENT_CELL(I) <= CURRENT_CELL(I-1);
        END LOOP;
        CURRENT_CELL(0) <= NEIGHBORHOOD_CELL(9, 9);
        ------------------------------------------------------------
		
		-- BINARY ADDER TREE FOR TOTAL STATES SUM ------------------
		FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 0 LOOP
			-- LOOP FOR EACH COLUMN:
			FOR I IN (NEIGHBORHOOD_SIZE-1)/2 DOWNTO 1 LOOP -- 19 = 2*9 + 1, 9 SUM RESULTS
				SUM_LAYER_0(I, J) <= NEIGHBORHOOD_REPLICA(2*I, J) + NEIGHBORHOOD_REPLICA(2*I-1, J);
			END LOOP;
			
			SUM_LAYER_0(0, J) <= NEIGHBORHOOD_REPLICA(0, J); 
			
			FOR I IN 4 DOWNTO 0 LOOP 
				SUM_LAYER_1(I, J) <= SUM_LAYER_0(2*I+1, J) + SUM_LAYER_0(2*I, J);
			END LOOP;
			
			SUM_LAYER_2(2, J) <= SUM_LAYER_1(4, J) + SUM_LAYER_1(3, J);
			SUM_LAYER_2(1, J) <= SUM_LAYER_1(2, J) + SUM_LAYER_1(1, J);
			SUM_LAYER_2(0, J) <= SUM_LAYER_1(0, J);
			
			SUM_LAYER_3(1, J) <= SUM_LAYER_2(2, J) + SUM_LAYER_2(1, J);
			SUM_LAYER_3(0, J) <= SUM_LAYER_2(0, J);
			
			SUM(J) <= SUM_LAYER_3(1, J) + SUM_LAYER_3(0, J);
		END LOOP;
		
		-- SUM(J) CONTAINS THE SUM OF COLUMN J
		-- ADDER TREE FOR THE SUM OF EACH COLUMN:
		FOR I IN (NEIGHBORHOOD_SIZE-1)/2 DOWNTO 1 LOOP 
			COLUMN_SUM_LAYER_0(I) <= SUM(2*I) + SUM(2*I-1);
		END LOOP;
		COLUMN_SUM_LAYER_0(0) <= SUM(0); 
		
		FOR I IN 4 DOWNTO 0 LOOP 
			COLUMN_SUM_LAYER_1(I) <= COLUMN_SUM_LAYER_0(2*I+1) + COLUMN_SUM_LAYER_0(2*I);
		END LOOP;
		
		COLUMN_SUM_LAYER_2(2) <= COLUMN_SUM_LAYER_1(4) + COLUMN_SUM_LAYER_1(3);
		COLUMN_SUM_LAYER_2(1) <= COLUMN_SUM_LAYER_1(2) + COLUMN_SUM_LAYER_1(1);
		COLUMN_SUM_LAYER_2(0) <= COLUMN_SUM_LAYER_1(0);
		
		COLUMN_SUM_LAYER_3(1) <= COLUMN_SUM_LAYER_2(2) + COLUMN_SUM_LAYER_2(1);
		COLUMN_SUM_LAYER_3(0) <= COLUMN_SUM_LAYER_2(0);
		
		TOTAL_SUM <= COLUMN_SUM_LAYER_3(1) + COLUMN_SUM_LAYER_3(0);
		------------------------------------------------------------
		
		-- BINARY ADDER TREE FOR TOTAL INFECTED CELLS SUM ------------------
		FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 0 LOOP
			-- LOOP FOR EACH COLUMN:
			FOR I IN (NEIGHBORHOOD_SIZE-1)/2 DOWNTO 1 LOOP -- 19 = 2*9 + 1, 9 SUM RESULTS
				INFECTED_SUM_LAYER_0(I, J) <= INFECTED_CELL(2*I, J) + INFECTED_CELL(2*I-1, J);
			END LOOP;
			
			INFECTED_SUM_LAYER_0(0, J) <= INFECTED_CELL(0, J); 
			
			FOR I IN 4 DOWNTO 0 LOOP 
				INFECTED_SUM_LAYER_1(I, J) <= INFECTED_SUM_LAYER_0(2*I+1, J) + INFECTED_SUM_LAYER_0(2*I, J);
			END LOOP;
			
			INFECTED_SUM_LAYER_2(2, J) <= INFECTED_SUM_LAYER_1(4, J) + INFECTED_SUM_LAYER_1(3, J);
			INFECTED_SUM_LAYER_2(1, J) <= INFECTED_SUM_LAYER_1(2, J) + INFECTED_SUM_LAYER_1(1, J);
			INFECTED_SUM_LAYER_2(0, J) <= INFECTED_SUM_LAYER_1(0, J);
			
			INFECTED_SUM_LAYER_3(1, J) <= INFECTED_SUM_LAYER_2(2, J) + INFECTED_SUM_LAYER_2(1, J);
			INFECTED_SUM_LAYER_3(0, J) <= INFECTED_SUM_LAYER_2(0, J);
			
			INFECTED_SUM(J) <= INFECTED_SUM_LAYER_3(1, J) + INFECTED_SUM_LAYER_3(0, J);
		END LOOP;
		
		-- SUM(J) CONTAINS THE SUM OF COLUMN J
		-- ADDER TREE FOR THE SUM OF EACH COLUMN:
		FOR I IN (NEIGHBORHOOD_SIZE-1)/2 DOWNTO 1 LOOP 
			INFECTED_COLUMN_SUM_LAYER_0(I) <= INFECTED_SUM(2*I) + INFECTED_SUM(2*I-1);
		END LOOP;
		
		INFECTED_COLUMN_SUM_LAYER_0(0) <= INFECTED_SUM(0); 
		
		FOR I IN 4 DOWNTO 0 LOOP 
			INFECTED_COLUMN_SUM_LAYER_1(I) <= INFECTED_COLUMN_SUM_LAYER_0(2*I+1) + INFECTED_COLUMN_SUM_LAYER_0(2*I);
		END LOOP;
		
		INFECTED_COLUMN_SUM_LAYER_2(2) <= INFECTED_COLUMN_SUM_LAYER_1(4) + INFECTED_COLUMN_SUM_LAYER_1(3);
		INFECTED_COLUMN_SUM_LAYER_2(1) <= INFECTED_COLUMN_SUM_LAYER_1(2) + INFECTED_COLUMN_SUM_LAYER_1(1);
		INFECTED_COLUMN_SUM_LAYER_2(0) <= INFECTED_COLUMN_SUM_LAYER_1(0);
		
		INFECTED_COLUMN_SUM_LAYER_3(1) <= INFECTED_COLUMN_SUM_LAYER_2(2) + INFECTED_COLUMN_SUM_LAYER_2(1);
		INFECTED_COLUMN_SUM_LAYER_3(0) <= INFECTED_COLUMN_SUM_LAYER_2(0);
		
		INFECTED_TOTAL_SUM <= INFECTED_COLUMN_SUM_LAYER_3(1) + INFECTED_COLUMN_SUM_LAYER_3(0);
		------------------------------------------------------------
		
		-- STATE TRANSITION RULE -----------------------------------
		IF CURRENT_CELL(10) = 0 then
		    IF INFECTED_TOTAL_SUM/64 > 255 THEN
		        DATA_OUT <= (OTHERS => '1'); -- 255
		    ELSE
		        DATA_OUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(INFECTED_TOTAL_SUM/64, 8));
		    END IF;
		ELSIF CURRENT_CELL(10) = 255 THEN 
			DATA_OUT <= (OTHERS => '0');
		ELSE
		    IF TOTAL_SUM/1024+5 > 255 THEN    
		        DATA_OUT <= (OTHERS => '1'); -- 255
		    ELSE 
		        DATA_OUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(TOTAL_SUM/1024+5, 8));
		    END IF;
		END IF;
		------------------------------------------------------------
		
		FOR I IN ((NEIGHBORHOOD_SIZE-1)/2)+12 DOWNTO 1 LOOP
            DATA_VALID_SIGNAL(I) <= DATA_VALID_SIGNAL(I-1);
        END LOOP;
        DATA_VALID_SIGNAL(0) <= READ_EN;		
		
	END PROCESS;
		
	DATA_OUT_VALID <= DATA_VALID_SIGNAL(((NEIGHBORHOOD_SIZE-1)/2)+12);	
		------------------------------------------------------------
	
END BEHAVIORAL;
	