----------------------------------------------------------------------------------
-- TECHNICAL UNIVERSITY OF CRETE
-- NICK KYPARISSAS
--
-- CREATE DATE: JUNE 2018
-- MODULE: GRAPHICS_CTRL 
-- PROJECT NAME: A Parallel Framework for Simulating Cellular Automata on FPGA Logic
-- XILINX OPEN HARDWARE 2018 ENTRY
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY GRAPHICS_CTRL IS
    GENERIC (
        COLOR_BITS : INTEGER := 4
    );    
	PORT ( 
		CLK 		: IN STD_LOGIC; -- @ 148.5 MHZ
		RST 		: IN STD_LOGIC;
		HS          : OUT STD_LOGIC;
        VS          : OUT STD_LOGIC;
        R           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        G           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        B           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		MEM_DATA	: IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		MEM_EN		: OUT STD_LOGIC;
		MEM_ACCESS_REQUEST : OUT STD_LOGIC;
		NEW_FRAME_LINE_REQUEST : OUT STD_LOGIC
	);
END GRAPHICS_CTRL;

ARCHITECTURE BEHAVIORAL OF GRAPHICS_CTRL IS
	--SIGNALS
	TYPE STD_LOGIC_ARRAY_2X12 IS ARRAY (2 DOWNTO 0) OF STD_LOGIC_VECTOR(11 DOWNTO 0); 
    SIGNAL HCWX_SIGNAL : STD_LOGIC_ARRAY_2X12;
    TYPE STD_LOGIC_ARRAY_2X11 IS ARRAY (2 DOWNTO 0) OF STD_LOGIC_VECTOR(10 DOWNTO 0); 
    SIGNAL VCWX_SIGNAL          : STD_LOGIC_ARRAY_2X11;
    SIGNAL HS_SIGNAL, VS_SIGNAL : STD_LOGIC_VECTOR(1 DOWNTO 0);
	
	BEGIN
	
	FHD_COLOR_CONTROLLER : ENTITY WORK.FHD_COLOR_CTRL
	    GENERIC MAP( 
	       COLOR_BITS => COLOR_BITS 
	    )
		PORT MAP(
			RST => RST,
			CLK => CLK,
			HCOUNT => HCWX_SIGNAL(2),
			VCOUNT => VCWX_SIGNAL(2),
			MEM_DATA => MEM_DATA,
			MEM_EN => MEM_EN, 
			RED => R,
			GREEN => G,
			BLUE => B
		);

	FHD_SYNC_CONTROLLER :  ENTITY WORK.FHD_CTRL
		PORT MAP(
			RST => RST, 
			CLK => CLK,
			HS => HS_SIGNAL(0),
			VS => VS_SIGNAL(0),
			HCOUNT => HCWX_SIGNAL(0),
			VCOUNT => VCWX_SIGNAL(0)    
		);
	
	PROCESS 
	BEGIN
		
		WAIT UNTIL RISING_EDGE(CLK);			
		
		--- WE NEED PIPELINING TO REACH 148.5 MHz 
		HS <= HS_SIGNAL(1);
		HS_SIGNAL(1) <= HS_SIGNAL(0);
		--
		VS <= VS_SIGNAL(1);
		VS_SIGNAL(1) <= VS_SIGNAL(0);
		--
		HCWX_SIGNAL(2) <= HCWX_SIGNAL(1);
		HCWX_SIGNAL(1) <= HCWX_SIGNAL(0);
		--
		VCWX_SIGNAL(2) <= VCWX_SIGNAL(1);
		VCWX_SIGNAL(1) <= VCWX_SIGNAL(0);
		-- 
		
		IF UNSIGNED(HCWX_SIGNAL(1)) > 1700 AND UNSIGNED(VCWX_SIGNAL(1)) = 1125 THEN
		  NEW_FRAME_LINE_REQUEST <= '1'; 
		ELSE
		  NEW_FRAME_LINE_REQUEST <= '0';
		END IF; 
		
		IF UNSIGNED(HCWX_SIGNAL(1)) > 1700 AND (UNSIGNED(VCWX_SIGNAL(1)) < 1079 OR UNSIGNED(VCWX_SIGNAL(1)) = 1125) THEN
            MEM_ACCESS_REQUEST <= '1';
        ELSE
            MEM_ACCESS_REQUEST <= '0';
        END IF;    
        
	END PROCESS;
	
END BEHAVIORAL;