----------------------------------------------------------------------------------
-- TECHNICAL UNIVERSITY OF CRETE
-- NICK KYPARISSAS
--
-- CREATE DATE: JUNE 2018
-- MODULE: GRID LINES BUFFER
-- PROJECT NAME: A Parallel Framework for Simulating Cellular Automata on FPGA Logic
-- XILINX OPEN HARDWARE 2018 ENTRY
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY GRID_LINES_BUFFER IS
	GENERIC (
        CELL_SIZE  			: INTEGER := 4;		
		BURST_SIZE 			: INTEGER := 128;
		GRID_X				: INTEGER := 1920;
		GRID_Y				: INTEGER := 1080;
		NUMBER_OF_BURSTS_PER_LINE 	: INTEGER := 60; -- GRID_X * CELL_SIZE / BURST_SIZE;
        NEIGHBORHOOD_SIZE  	: INTEGER := 5); 
    PORT (
        CLK_200        	: IN STD_LOGIC; -- SYSTEM CLOCK
		UI_CLK        	: IN STD_LOGIC; -- SYSTEM CLOCK
		RST         	: IN STD_LOGIC; -- HIGH ACTIVE SYNCHRONOUS RESET
		WRITE_EN		: IN STD_LOGIC;
        DATA_IN     	: IN STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0);
        MEMORY_ACCESS_GRANTED : IN STD_LOGIC;
        DATA_OUT   		: OUT STD_LOGIC_VECTOR((NEIGHBORHOOD_SIZE*CELL_SIZE)-1 DOWNTO 0);
        DATA_OUT_VALID 	: OUT STD_LOGIC -- WHEN DATA_OUT_VALID = 1, THE ARRAY IS BEING DRAINED, ONE DATA_OUT COLUMN PER CLK CYCLE
        ); 
END GRID_LINES_BUFFER;

ARCHITECTURE BEHAVIORAL OF GRID_LINES_BUFFER IS
	
	SIGNAL WRITE_ADDRESS_COUNTER : INTEGER RANGE 0 TO NUMBER_OF_BURSTS_PER_LINE-1 := 0;
	SIGNAL READ_ADDRESS_COUNTER : INTEGER RANGE 0 TO GRID_X-1 := 0;
	
	TYPE CRAPPY_SIGNAL IS ARRAY (NEIGHBORHOOD_SIZE DOWNTO 0) OF STD_LOGIC_VECTOR(0 DOWNTO 0); 
	SIGNAL WRITE_ENABLE : CRAPPY_SIGNAL;
	
	SIGNAL WRITE_ADDRESS : STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL READ_ADDRESS : STD_LOGIC_VECTOR(10 DOWNTO 0);
	
	TYPE INTEGER_SYNCHRONIZER_1 IS ARRAY (1 DOWNTO 0) OF INTEGER RANGE 0 TO GRID_Y;
	SIGNAL TOTAL_NUM_OF_FILLED_LINES : INTEGER_SYNCHRONIZER_1;
	
	SIGNAL DATA_OUT_VALID_SIGNAL : STD_LOGIC_VECTOR(NEIGHBORHOOD_SIZE-1 DOWNTO 0) := (OTHERS => '0');
	
	TYPE INTEGER_SYNCHRONIZER_2 IS ARRAY (1 DOWNTO 0) OF INTEGER RANGE 0 TO NEIGHBORHOOD_SIZE;
	SIGNAL LINE_BEING_FILLED	: INTEGER_SYNCHRONIZER_2;
	
	TYPE STD_LOGIC_ARRAY IS ARRAY (NEIGHBORHOOD_SIZE-1 DOWNTO 0, NEIGHBORHOOD_SIZE DOWNTO 0) OF STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
	SIGNAL LINE_DATA : STD_LOGIC_ARRAY; 
	
	TYPE INTEGER_ARRAY IS ARRAY (NEIGHBORHOOD_SIZE-1 DOWNTO 0, NEIGHBORHOOD_SIZE-1 DOWNTO 0) OF INTEGER RANGE 0 TO NEIGHBORHOOD_SIZE;
	SIGNAL LINES_BEING_DRAINED : INTEGER_ARRAY;
	
	SIGNAL SYNC_CONTROL : STD_LOGIC := '0';
	
	TYPE STATE IS (RESET, WAIT_FOR_BUFFER_FILL, BUFFER_DRAIN);
	SIGNAL FSM_STATE : STATE;	
	
	COMPONENT LINE_BUFFER_4b 
  	PORT (
	    clka : IN STD_LOGIC;
	    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
	    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	    dina : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
	    clkb : IN STD_LOGIC;
	    addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
	    doutb : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  	);
	END COMPONENT;
	
	COMPONENT LINE_BUFFER_8B 
    PORT (
        clka : IN STD_LOGIC;
        wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
        addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
        dina : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
        clkb : IN STD_LOGIC;
        addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
        doutb : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
      );
    END COMPONENT;

BEGIN
	
	GENERATE_LINE_BUFFERS: for I in 0 to NEIGHBORHOOD_SIZE generate 
	-- 0 to NEIGHBORHOOD_SIZE-1 LINES + ONE FOR BUFFERING
		LINE_BUFFER_4:	IF (CELL_SIZE = 4) GENERATE
            LINE_BUFFER: LINE_BUFFER_4b 
            PORT MAP(
                clka => UI_CLK,
                wea => WRITE_ENABLE(I),
                addra => WRITE_ADDRESS(5 DOWNTO 0),
                dina => DATA_IN,
                clkb => CLK_200,
                addrb => READ_ADDRESS,
                doutb => LINE_DATA(0, I)
            ); 
  		END GENERATE LINE_BUFFER_4;
  		
  		LINE_BUFFER_8:	IF (CELL_SIZE = 8) GENERATE
            LINE_BUFFER: LINE_BUFFER_8b 
            PORT MAP(
                clka => UI_CLK,
                wea => WRITE_ENABLE(I),
                addra => WRITE_ADDRESS,
                dina => DATA_IN,
                clkb => CLK_200,
                addrb => READ_ADDRESS,
                doutb => LINE_DATA(0, I)
            );
        END GENERATE LINE_BUFFER_8;
	end generate GENERATE_LINE_BUFFERS;
	
	SYNCHRONIZER: ENTITY WORK.SYNCHRONIZER
	GENERIC MAP (
		GRID_Y => GRID_Y,
        NEIGHBORHOOD_SIZE => NEIGHBORHOOD_SIZE
    ) 
	PORT MAP (
		CLK_RX => CLK_200,
		RST => RST,
		--
		CONTROL => SYNC_CONTROL,
		DATA_IN_1 => TOTAL_NUM_OF_FILLED_LINES(0),
		DATA_OUT_1 => TOTAL_NUM_OF_FILLED_LINES(1),
		-- SYNCHRONIZING COMMUNICATING FSM SIGNALS:
		DATA_IN_2 => LINE_BEING_FILLED(0),
		DATA_OUT_2 => LINE_BEING_FILLED(1)
	);
	
	WRITE_ADDRESS <= STD_LOGIC_VECTOR(TO_UNSIGNED(WRITE_ADDRESS_COUNTER, WRITE_ADDRESS'LENGTH));
    READ_ADDRESS <= STD_LOGIC_VECTOR(TO_UNSIGNED(READ_ADDRESS_COUNTER, READ_ADDRESS'LENGTH));
    
	WRITE: PROCESS
	BEGIN
		
		WAIT UNTIL RISING_EDGE(UI_CLK);		
		
		IF RST = '1' THEN
			WRITE_ADDRESS_COUNTER <= 0;
			LINE_BEING_FILLED(0) <= 0;
			TOTAL_NUM_OF_FILLED_LINES(0) <= 0;
			SYNC_CONTROL <= '0';
		ELSE
			IF WRITE_EN = '1' AND MEMORY_ACCESS_GRANTED = '1' THEN
				IF WRITE_ADDRESS_COUNTER = NUMBER_OF_BURSTS_PER_LINE-1 THEN
					WRITE_ADDRESS_COUNTER <= 0;
					IF LINE_BEING_FILLED(0) = NEIGHBORHOOD_SIZE THEN 
					-- SOME SYNTHESIZERS WOULD CALCULATE THE OVERFLOW, BUT WE CHOOSE TO BE EXPLICIT
						LINE_BEING_FILLED(0) <= 0;
					ELSE
						LINE_BEING_FILLED(0) <= LINE_BEING_FILLED(0) + 1;
					END IF;
					-- NOTIFYING THE READER THERE IS A NEW LINE_BEING_FILLED VALUE
					TOTAL_NUM_OF_FILLED_LINES(0) <= TOTAL_NUM_OF_FILLED_LINES(0) + 1;
					SYNC_CONTROL <= '1';
				ELSE
					WRITE_ADDRESS_COUNTER <= WRITE_ADDRESS_COUNTER + 1;
					SYNC_CONTROL <= '0';
				END IF;
			ELSIF MEMORY_ACCESS_GRANTED = '0' AND TOTAL_NUM_OF_FILLED_LINES(0) = GRID_Y THEN
			    -- NO ISSUE WITH COMMUNICATING WITH THE READING PROCESS:
			    -- LINE_BEING_FILLED(0) <= 0; AFTER THAT PROCESS HAS STARTED DRAINING THE BUFFER
			    TOTAL_NUM_OF_FILLED_LINES(0) <= 0;
			    LINE_BEING_FILLED(0) <= 0;
			    SYNC_CONTROL <= '1';
			ELSE 
				WRITE_ADDRESS_COUNTER <= WRITE_ADDRESS_COUNTER;
				TOTAL_NUM_OF_FILLED_LINES(0) <= TOTAL_NUM_OF_FILLED_LINES(0);
				LINE_BEING_FILLED(0) <= LINE_BEING_FILLED(0);
				SYNC_CONTROL <= '0';
			END IF;
		END IF;
	
	END PROCESS WRITE;
	
	SETTING_WREN: PROCESS(WRITE_EN, LINE_BEING_FILLED(0))
	BEGIN
		for I in 0 to NEIGHBORHOOD_SIZE LOOP
			IF I = LINE_BEING_FILLED(0) THEN
				WRITE_ENABLE(I)(0) <= WRITE_EN;
			ELSE
				WRITE_ENABLE(I)(0) <= '0';
			END IF;
		END LOOP;
	END PROCESS SETTING_WREN;
	
	READ: PROCESS
	BEGIN
		
		WAIT UNTIL RISING_EDGE(CLK_200);
		
		IF RST = '1' THEN
			FSM_STATE <= RESET;
		ELSE
			CASE FSM_STATE IS 
			WHEN RESET =>
				FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
					LINES_BEING_DRAINED(0, I) <= I;
				END LOOP;
				READ_ADDRESS_COUNTER <= 0;
				DATA_OUT_VALID <= '0';
				DATA_OUT_VALID_SIGNAL <= (OTHERS => '0');
				-- TEST
				--TOTAL_NUM_OF_DRAINED_LINES <= 0;
				FSM_STATE <= WAIT_FOR_BUFFER_FILL;
			WHEN WAIT_FOR_BUFFER_FILL =>
				IF TOTAL_NUM_OF_FILLED_LINES(1) >= NEIGHBORHOOD_SIZE AND LINES_BEING_DRAINED(0, NEIGHBORHOOD_SIZE-1) /= LINE_BEING_FILLED(1) THEN --AND TOTAL_NUM_OF_DRAINED_LINES /= (GRID_Y)-(NEIGHBORHOOD_SIZE-1) THEN 
					-- IF THERE ARE ENOUGH LINES IN THE BUFFER 
					-- AND THE LINE WE ARE ABOUT TO DRAIN IS NOT THE ONE THAT'S BEING FILLED
					-- AND A NEW FRAME HAS BEING LOADED
					FSM_STATE <= BUFFER_DRAIN;
				ELSE
					FSM_STATE <= FSM_STATE;  
				END IF;
				
				-- NEW FRAME: RESETTING WHICH LINES TO DRAIN
                IF TOTAL_NUM_OF_FILLED_LINES(1) = 0 THEN
                    FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
                       LINES_BEING_DRAINED(0, I) <= I;
                    END LOOP; 
                END IF;
				
				DATA_OUT_VALID_SIGNAL(0) <= '0';

			WHEN BUFFER_DRAIN =>				
				
				IF READ_ADDRESS_COUNTER = GRID_X-1 THEN
					READ_ADDRESS_COUNTER <= 0;
					FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
						-- MOST SYNTHESIZERS WOULD CALCULATE THE OVERFLOW, BUT WE CHOOSE TO BE EXPLICIT
						IF LINES_BEING_DRAINED(0, I) = NEIGHBORHOOD_SIZE THEN
							LINES_BEING_DRAINED(0, I) <= 0;
						ELSE
							LINES_BEING_DRAINED(0, I) <= LINES_BEING_DRAINED(0, I) + 1;
						END IF;
					END LOOP;				
					FSM_STATE <= WAIT_FOR_BUFFER_FILL;  
                
				ELSE
					READ_ADDRESS_COUNTER <= READ_ADDRESS_COUNTER + 1;
					DATA_OUT_VALID_SIGNAL(0) <= '1';
					FSM_STATE <= FSM_STATE;
				END IF;
                                    
			END CASE;
		END IF;
		
		-- PIPELINING REGISTERS FOR THE OUTPUTS
		-- AS THE SIZE OF NEIGHBORHOOD RISES, THE NUMBER OF BRAM MODULES RISES AS WELL
		-- ROUTING NEEDS MORE SLACK
		DATA_OUT_VALID <= DATA_OUT_VALID_SIGNAL(NEIGHBORHOOD_SIZE-1);
		FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 1 LOOP	
			DATA_OUT_VALID_SIGNAL(J) <= DATA_OUT_VALID_SIGNAL(J-1);
	    END LOOP;
		-- THE LINES BEING DRAINED CHANGE OVER TIME: (0, LINES_BEING_DRAINED(I))
        
        FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP	
            DATA_OUT(((I+1)*CELL_SIZE)-1 DOWNTO (I*CELL_SIZE)) <= LINE_DATA(NEIGHBORHOOD_SIZE-1,  LINES_BEING_DRAINED(NEIGHBORHOOD_SIZE-1, I)); 
        END LOOP;
        
		L_1: FOR I IN 0 TO NEIGHBORHOOD_SIZE LOOP
		    L_2: FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 1 LOOP	
                LINE_DATA(J, I) <= LINE_DATA(J-1, I);
            END LOOP L_2;
        END LOOP L_1;
        
        L_3: FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
        	L_4: FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 1 LOOP	
        		LINES_BEING_DRAINED(J, I) <= LINES_BEING_DRAINED(J-1, I);
        	END LOOP L_4;
        END LOOP L_3;

	END PROCESS READ;
	
END BEHAVIORAL;