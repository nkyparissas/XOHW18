----------------------------------------------------------------------------------
-- TECHNICAL UNIVERSITY OF CRETE
-- NICK KYPARISSAS
--
-- CREATE DATE: JUNE 2018
-- MODULE: MEMORY ACCESS ARBITRATOR
-- PROJECT NAME: A Parallel Framework for Simulating Cellular Automata on FPGA Logic
-- XILINX OPEN HARDWARE 2018 ENTRY
----------------------------------------------------------------------------------

-----------------------------------------------------------------------------
-- NOT THAT EACH STATE CHANGES ONLY IT'S OWN MUX_SEL 
-- WE NEED A CYCLE DELAY BETWEEN ACCESS GRANTED AND MUX FOR TAGGING
-----------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MEMORY_ACCESS_ARBITRATOR IS
    PORT ( 	CLK						: IN STD_LOGIC;	-- UI CLOCK 
			RST 					: IN STD_LOGIC;
			-- INIT SIGNALS --
			INIT_COMPLETE			: IN STD_LOGIC;
			-- GRAPHICS SIGNALS	--
			GRAPHICS_REQ			: IN STD_LOGIC;
			GRAPHICS_NEW_FRAME_REQ	: IN STD_LOGIC;
			GRAPHICS_ACCESS_GRANTED	: OUT STD_LOGIC;
			-- DATAPATH WRITE SIGNALS --
			WRITE_BACK_ACCESS_GRANTED	: OUT STD_LOGIC;
			-- DDR SIGNALS --
			APP_CMD_SELECT 		: OUT STD_LOGIC_VECTOR(1 DOWNTO 0); -- 00: INIT, 01: GRAPHICS AND LINES BUFFER, 10: DATAPATH WRITE
			APP_WRITE_SELECT		: OUT STD_LOGIC--; -- 0: INIT, 1: WRITING BUFFER

	);
END MEMORY_ACCESS_ARBITRATOR;

ARCHITECTURE BEHAVIORAL OF MEMORY_ACCESS_ARBITRATOR IS
	
    SIGNAL GRAPHICS_REQ_SIGNAL, GRAPHICS_NEW_FRAME_REQ_SIGNAL : STD_LOGIC_VECTOR(1 DOWNTO 0);
	TYPE STATE IS (RESET, WAIT_FOR_FRAME_ALIGNMENT, GRAPHICS_AND_LINES_BUFFER, WRITE_BACK);
		SIGNAL FSM_STATE : STATE;

BEGIN
    
	-- THE FOLLOWING FSM HANDLES THE DATA BEING RECEIVED  
	DATA_IN_FLOW_CONTROL: PROCESS 
		BEGIN
		
		WAIT UNTIL CLK'EVENT AND CLK = '1';
		
		IF (RST = '1') THEN  
			FSM_STATE <= RESET;    
		ELSE
			CASE FSM_STATE IS 
			WHEN RESET => 
				GRAPHICS_ACCESS_GRANTED	<= '0';
				WRITE_BACK_ACCESS_GRANTED <= '0';
				-- DDR SIGNALS --
				APP_CMD_SELECT <= "00";
				APP_WRITE_SELECT <= '0';

				FSM_STATE <= WAIT_FOR_FRAME_ALIGNMENT;
			WHEN WAIT_FOR_FRAME_ALIGNMENT =>
				IF (GRAPHICS_NEW_FRAME_REQ_SIGNAL(0) = '1' AND INIT_COMPLETE = '1') THEN 
				-- WE HAVE TO MAKE SURE THAT THE FIRST LINE OF THE BUFFER WILL BE LOADED IN OUR GRAPHICS BUFFER BEFORE ANY OTHER LINE
					FSM_STATE <= GRAPHICS_AND_LINES_BUFFER;
					APP_WRITE_SELECT <= '1';
				ELSE 
					FSM_STATE <= WAIT_FOR_FRAME_ALIGNMENT;
				END IF;
			WHEN GRAPHICS_AND_LINES_BUFFER =>
				IF (GRAPHICS_REQ_SIGNAL(0) = '1' OR GRAPHICS_NEW_FRAME_REQ_SIGNAL(0) = '1') THEN
                    WRITE_BACK_ACCESS_GRANTED    <= '0';
                    GRAPHICS_ACCESS_GRANTED    <= '1';
					APP_CMD_SELECT <= "01"; -- GRAPHICS AND LINES BUFFER
					FSM_STATE <= FSM_STATE;
				ELSE
                    WRITE_BACK_ACCESS_GRANTED    <= '0'; 
                    GRAPHICS_ACCESS_GRANTED    <= '0';
                    FSM_STATE <= WRITE_BACK;
				END IF;  				
			WHEN WRITE_BACK =>	
				IF (GRAPHICS_REQ_SIGNAL(0) = '1' OR GRAPHICS_NEW_FRAME_REQ_SIGNAL(0) = '1') THEN
                    WRITE_BACK_ACCESS_GRANTED    <= '0';
                    GRAPHICS_ACCESS_GRANTED    <= '0';
					FSM_STATE <= GRAPHICS_AND_LINES_BUFFER;
				ELSE
                    WRITE_BACK_ACCESS_GRANTED    <= '1'; 
                    GRAPHICS_ACCESS_GRANTED    <= '0';
					APP_CMD_SELECT <= "10"; -- WRITE_BACK  
					FSM_STATE <= FSM_STATE;
				END IF;
			END CASE;
		END IF;
	END PROCESS DATA_IN_FLOW_CONTROL;
	
	-- GRAPHICS CONTROLLER OPERATES IN A DIFFERENT CLOCK DOMAIN
	GRAPHICS_AND_DDR_ACCESS_CONTROL_SYNCHRONIZATION: PROCESS 
	BEGIN
	
		WAIT UNTIL CLK'EVENT AND CLK = '1';
		
		IF (RST = '1') THEN
			GRAPHICS_REQ_SIGNAL <= (OTHERS => '0');
			GRAPHICS_NEW_FRAME_REQ_SIGNAL <= (OTHERS => '0');
		ELSE
			GRAPHICS_REQ_SIGNAL(0) <= GRAPHICS_REQ_SIGNAL(1);
			GRAPHICS_REQ_SIGNAL(1) <= GRAPHICS_REQ;
			GRAPHICS_NEW_FRAME_REQ_SIGNAL(0) <= GRAPHICS_NEW_FRAME_REQ_SIGNAL(1);
			GRAPHICS_NEW_FRAME_REQ_SIGNAL(1) <= GRAPHICS_NEW_FRAME_REQ;
		END IF;		
	END PROCESS GRAPHICS_AND_DDR_ACCESS_CONTROL_SYNCHRONIZATION;
	
END BEHAVIORAL;